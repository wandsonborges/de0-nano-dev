rodrigo@thomson.7111477660155