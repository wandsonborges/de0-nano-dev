rodrigo@debian.2917:1553254025