module burst_read_wf
  (
   clk,
   reset,

   master_address,
   master_read,
   master_readdata,
   master_burstcount,
   //master_byteenable,
   master_waitrequest,
   master_readdatavalid,

   ctrl_start,
   ctrl_baseaddress,
   ctrl_burstcount,
   ctrl_busy,
   ctrl_readdatavalid,
   ctrl_readdata
   );


  parameter ADDRESS_WIDTH = 32;          // derived parameter (using system info)
  parameter LENGTH_WIDTH = 32;           // any value from 4-32 (larger the value the slower the logic will be), LENGTH_WIDTH shouldn't be larger than ADDRESS_WIDTH and should be reduced to increase the Fmax of the master.
  parameter DATA_WIDTH = 32;             // 16, 32, 64, 128, 256, 512, 1024 are valid choices
  parameter BYTE_ENABLE_WIDTH = 4;       // derived parameter
  parameter BYTE_ENABLE_WIDTH_LOG2 = 2;  // derived parameter
  parameter BURST_COUNT = 2;         // must be a multiple of 2 between 2 and 1024, when bursting is disabled this value must be set to 1
  parameter BURST_WIDTH = 2;             // derived parameter


   localparam ST_START = 3'b001, ST_WAITREQUEST = 3'b010, ST_BURST = 3'b100;
   
   input clk;
   input reset;					// 

   
   output reg [ADDRESS_WIDTH-1:0] master_address;
   output reg master_read;
   //output reg 				   master_beginbursttransfer;
   output reg [BURST_WIDTH-1:0] master_burstcount;
   //output wire [BYTE_ENABLE_WIDTH-1:0] master_byteenable;
   input 	   master_waitrequest;
   input 	   master_readdatavalid;
   input [DATA_WIDTH-1:0] master_readdata;
	   

   input 	   ctrl_start;
   input [ADDRESS_WIDTH-1:0] 	   ctrl_baseaddress;
   input [BURST_WIDTH-1:0] 		   ctrl_burstcount;
   output reg  ctrl_busy;
   output wire ctrl_readdatavalid;
   output wire [DATA_WIDTH-1:0] ctrl_readdata;
   



   reg [BURST_WIDTH-1:0] burstCount;
   reg [2:0] 			 state;
   

   wire 				 local_ctrl_start;
   


   assign local_ctrl_start = ~ctrl_busy;
   
   // always @(ctrl_busy)
   // 	 begin
   // 		if (ctrl_busy == 0)
   // 		  begin
   // 			 local_ctrl_start = 1;
   // 		  end


   
   

   always @(posedge clk or posedge reset)
	 begin
		if (reset == 1)
		  begin
				  master_address <= 0;
				  master_burstcount <= 0;
				  master_read <= 1'b0;
				  ctrl_busy <= 1'b0;
				  burstCount <= 0;
			 state <= ST_START;
			 
		  end
		else
		  begin
			 case (state)
			   ST_START:
				 if (local_ctrl_start == 1)
				   begin
					  master_address <= 32'h39000000;
 //ctrl_baseaddress;
					  master_burstcount <= 8;
 //ctrl_burstcount;
					  master_read <= 1'b1;

					  ctrl_busy <= 1'b1;

					  burstCount <= 0;
					  state <= ST_WAITREQUEST;
					  
				   end // if (local_ctrl_start == 1)
			   ST_WAITREQUEST:
				 if (master_waitrequest == 0)
				   begin
					  master_read <= 1'b0;
					  
					  state <= ST_BURST;
				   end
			   ST_BURST:
				 if (master_readdatavalid)
				   begin
					   //if (burstCount == (ctrl_burstcount-1))
					   if (burstCount == 7)
						 begin
							ctrl_busy <= 1'b0;
							burstCount <= 0;
							state <= ST_START;
							
						 end
					   else
						 begin
							burstCount <= burstCount + 1;
						 end
				   end // if (master_waitrequest == 0)
			   default:
				 state <= ST_START;
			   
			 endcase // case (state)
		  end
	 end		
					   
					   
   assign ctrl_readdatavalid = master_readdatavalid;
   assign ctrl_readdata = master_readdata;
   
   
				  
endmodule // burst_write_wf



   
