// cycloneV_soc.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module cycloneV_soc (
		input  wire        clk_clk,                         //                     clk.clk
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //                  hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                        .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                        .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                        .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                        .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                        .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                        .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                        .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                        .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                        .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                        .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                        .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                        .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                        .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                        .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                        .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                        .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                        .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                        .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                        .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                        .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                        .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                        .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                        .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                        .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                        .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                        .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                        .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                        .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                        .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                        .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                        .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                        .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                        .hps_io_uart0_inst_TX
		output wire [7:0]  led_external_connection_export,  // led_external_connection.export
		input  wire [7:0]  lwir_ul0304_datain,              //             lwir_ul0304.datain
		output wire        lwir_ul0304_syt,                 //                        .syt
		output wire        lwir_ul0304_syl,                 //                        .syl
		output wire        lwir_ul0304_syp,                 //                        .syp
		output wire [14:0] memory_mem_a,                    //                  memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                        .mem_ba
		output wire        memory_mem_ck,                   //                        .mem_ck
		output wire        memory_mem_ck_n,                 //                        .mem_ck_n
		output wire        memory_mem_cke,                  //                        .mem_cke
		output wire        memory_mem_cs_n,                 //                        .mem_cs_n
		output wire        memory_mem_ras_n,                //                        .mem_ras_n
		output wire        memory_mem_cas_n,                //                        .mem_cas_n
		output wire        memory_mem_we_n,                 //                        .mem_we_n
		output wire        memory_mem_reset_n,              //                        .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                        .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                        .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                        .mem_dqs_n
		output wire        memory_mem_odt,                  //                        .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                        .mem_dm
		input  wire        memory_oct_rzqin,                //                        .oct_rzqin
		input  wire        reset_reset_n,                   //                   reset.reset_n
		input  wire [3:0]  sw_external_connection_export,   //  sw_external_connection.export
		output wire        swir_v400_sensor_clk,            //               swir_v400.sensor_clk
		input  wire [7:0]  swir_v400_datain,                //                        .datain
		output wire        swir_v400_fsync,                 //                        .fsync
		output wire        swir_v400_lsync,                 //                        .lsync
		output wire        swir_v400_swir_pxl_clk_out       //                        .swir_pxl_clk_out
	);

	wire         pll_0_outclk0_clk;                                            // pll_0:outclk_0 -> [avalon_st_adapter_001:in_clk_0_clk, bridge_stSrcMmMaster_1:clk, mm_interconnect_4:pll_0_outclk0_clk, rst_controller_002:clk, swir_v400_0:pxl_clk_in]
	wire         pll_0_outclk1_clk;                                            // pll_0:outclk_1 -> [avalon_st_adapter:in_clk_0_clk, bridge_stSrcMmMaster_0:clk, lwir_ul0304_0:sensor_clk_in, mm_interconnect_4:pll_0_outclk1_clk, rst_controller_001:clk, swir_v400_0:sensor_clk_in]
	wire         bridge_stsrcmmmaster_1_avalon_master_waitrequest;             // mm_interconnect_0:bridge_stSrcMmMaster_1_avalon_master_waitrequest -> bridge_stSrcMmMaster_1:master_waitrequest
	wire  [31:0] bridge_stsrcmmmaster_1_avalon_master_address;                 // bridge_stSrcMmMaster_1:master_address -> mm_interconnect_0:bridge_stSrcMmMaster_1_avalon_master_address
	wire         bridge_stsrcmmmaster_1_avalon_master_write;                   // bridge_stSrcMmMaster_1:master_write -> mm_interconnect_0:bridge_stSrcMmMaster_1_avalon_master_write
	wire   [7:0] bridge_stsrcmmmaster_1_avalon_master_writedata;               // bridge_stSrcMmMaster_1:master_writedata -> mm_interconnect_0:bridge_stSrcMmMaster_1_avalon_master_writedata
	wire   [3:0] bridge_stsrcmmmaster_1_avalon_master_burstcount;              // bridge_stSrcMmMaster_1:master_burstcount -> mm_interconnect_0:bridge_stSrcMmMaster_1_avalon_master_burstcount
	wire         mm_interconnect_0_hps_0_f2h_sdram1_data_waitrequest;          // hps_0:f2h_sdram1_WAITREQUEST -> mm_interconnect_0:hps_0_f2h_sdram1_data_waitrequest
	wire  [29:0] mm_interconnect_0_hps_0_f2h_sdram1_data_address;              // mm_interconnect_0:hps_0_f2h_sdram1_data_address -> hps_0:f2h_sdram1_ADDRESS
	wire   [3:0] mm_interconnect_0_hps_0_f2h_sdram1_data_byteenable;           // mm_interconnect_0:hps_0_f2h_sdram1_data_byteenable -> hps_0:f2h_sdram1_BYTEENABLE
	wire         mm_interconnect_0_hps_0_f2h_sdram1_data_write;                // mm_interconnect_0:hps_0_f2h_sdram1_data_write -> hps_0:f2h_sdram1_WRITE
	wire  [31:0] mm_interconnect_0_hps_0_f2h_sdram1_data_writedata;            // mm_interconnect_0:hps_0_f2h_sdram1_data_writedata -> hps_0:f2h_sdram1_WRITEDATA
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram1_data_burstcount;           // mm_interconnect_0:hps_0_f2h_sdram1_data_burstcount -> hps_0:f2h_sdram1_BURSTCOUNT
	wire         bridge_stsrcmmmaster_0_avalon_master_waitrequest;             // mm_interconnect_1:bridge_stSrcMmMaster_0_avalon_master_waitrequest -> bridge_stSrcMmMaster_0:master_waitrequest
	wire  [31:0] bridge_stsrcmmmaster_0_avalon_master_address;                 // bridge_stSrcMmMaster_0:master_address -> mm_interconnect_1:bridge_stSrcMmMaster_0_avalon_master_address
	wire         bridge_stsrcmmmaster_0_avalon_master_write;                   // bridge_stSrcMmMaster_0:master_write -> mm_interconnect_1:bridge_stSrcMmMaster_0_avalon_master_write
	wire   [7:0] bridge_stsrcmmmaster_0_avalon_master_writedata;               // bridge_stSrcMmMaster_0:master_writedata -> mm_interconnect_1:bridge_stSrcMmMaster_0_avalon_master_writedata
	wire   [3:0] bridge_stsrcmmmaster_0_avalon_master_burstcount;              // bridge_stSrcMmMaster_0:master_burstcount -> mm_interconnect_1:bridge_stSrcMmMaster_0_avalon_master_burstcount
	wire         mm_interconnect_1_hps_0_f2h_sdram3_data_waitrequest;          // hps_0:f2h_sdram3_WAITREQUEST -> mm_interconnect_1:hps_0_f2h_sdram3_data_waitrequest
	wire  [29:0] mm_interconnect_1_hps_0_f2h_sdram3_data_address;              // mm_interconnect_1:hps_0_f2h_sdram3_data_address -> hps_0:f2h_sdram3_ADDRESS
	wire   [3:0] mm_interconnect_1_hps_0_f2h_sdram3_data_byteenable;           // mm_interconnect_1:hps_0_f2h_sdram3_data_byteenable -> hps_0:f2h_sdram3_BYTEENABLE
	wire         mm_interconnect_1_hps_0_f2h_sdram3_data_write;                // mm_interconnect_1:hps_0_f2h_sdram3_data_write -> hps_0:f2h_sdram3_WRITE
	wire  [31:0] mm_interconnect_1_hps_0_f2h_sdram3_data_writedata;            // mm_interconnect_1:hps_0_f2h_sdram3_data_writedata -> hps_0:f2h_sdram3_WRITEDATA
	wire   [7:0] mm_interconnect_1_hps_0_f2h_sdram3_data_burstcount;           // mm_interconnect_1:hps_0_f2h_sdram3_data_burstcount -> hps_0:f2h_sdram3_BURSTCOUNT
	wire  [31:0] addvector_0_avalon_rd1_1_1_1_readdata;                        // mm_interconnect_2:addVector_0_avalon_rd1_1_1_1_readdata -> addVector_0:masterrd1_readdata
	wire         addvector_0_avalon_rd1_1_1_1_waitrequest;                     // mm_interconnect_2:addVector_0_avalon_rd1_1_1_1_waitrequest -> addVector_0:masterrd1_waitrequest
	wire  [31:0] addvector_0_avalon_rd1_1_1_1_address;                         // addVector_0:masterrd1_address -> mm_interconnect_2:addVector_0_avalon_rd1_1_1_1_address
	wire         addvector_0_avalon_rd1_1_1_1_read;                            // addVector_0:masterrd1_read -> mm_interconnect_2:addVector_0_avalon_rd1_1_1_1_read
	wire         addvector_0_avalon_rd1_1_1_1_readdatavalid;                   // mm_interconnect_2:addVector_0_avalon_rd1_1_1_1_readdatavalid -> addVector_0:masterrd1_readdatavalid
	wire   [3:0] addvector_0_avalon_rd1_1_1_1_burstcount;                      // addVector_0:masterrd1_burstcount -> mm_interconnect_2:addVector_0_avalon_rd1_1_1_1_burstcount
	wire  [31:0] addvector_1_avalon_rd1_1_1_1_readdata;                        // mm_interconnect_2:addVector_1_avalon_rd1_1_1_1_readdata -> addVector_1:masterrd1_readdata
	wire         addvector_1_avalon_rd1_1_1_1_waitrequest;                     // mm_interconnect_2:addVector_1_avalon_rd1_1_1_1_waitrequest -> addVector_1:masterrd1_waitrequest
	wire  [31:0] addvector_1_avalon_rd1_1_1_1_address;                         // addVector_1:masterrd1_address -> mm_interconnect_2:addVector_1_avalon_rd1_1_1_1_address
	wire         addvector_1_avalon_rd1_1_1_1_read;                            // addVector_1:masterrd1_read -> mm_interconnect_2:addVector_1_avalon_rd1_1_1_1_read
	wire         addvector_1_avalon_rd1_1_1_1_readdatavalid;                   // mm_interconnect_2:addVector_1_avalon_rd1_1_1_1_readdatavalid -> addVector_1:masterrd1_readdatavalid
	wire   [3:0] addvector_1_avalon_rd1_1_1_1_burstcount;                      // addVector_1:masterrd1_burstcount -> mm_interconnect_2:addVector_1_avalon_rd1_1_1_1_burstcount
	wire  [31:0] addvector_0_avalon_rd2_readdata;                              // mm_interconnect_2:addVector_0_avalon_rd2_readdata -> addVector_0:masterrd2_readdata
	wire         addvector_0_avalon_rd2_waitrequest;                           // mm_interconnect_2:addVector_0_avalon_rd2_waitrequest -> addVector_0:masterrd2_waitrequest
	wire  [31:0] addvector_0_avalon_rd2_address;                               // addVector_0:masterrd2_address -> mm_interconnect_2:addVector_0_avalon_rd2_address
	wire         addvector_0_avalon_rd2_read;                                  // addVector_0:masterrd2_read -> mm_interconnect_2:addVector_0_avalon_rd2_read
	wire         addvector_0_avalon_rd2_readdatavalid;                         // mm_interconnect_2:addVector_0_avalon_rd2_readdatavalid -> addVector_0:masterrd2_readdatavalid
	wire   [3:0] addvector_0_avalon_rd2_burstcount;                            // addVector_0:masterrd2_burstcount -> mm_interconnect_2:addVector_0_avalon_rd2_burstcount
	wire  [31:0] addvector_1_avalon_rd2_readdata;                              // mm_interconnect_2:addVector_1_avalon_rd2_readdata -> addVector_1:masterrd2_readdata
	wire         addvector_1_avalon_rd2_waitrequest;                           // mm_interconnect_2:addVector_1_avalon_rd2_waitrequest -> addVector_1:masterrd2_waitrequest
	wire  [31:0] addvector_1_avalon_rd2_address;                               // addVector_1:masterrd2_address -> mm_interconnect_2:addVector_1_avalon_rd2_address
	wire         addvector_1_avalon_rd2_read;                                  // addVector_1:masterrd2_read -> mm_interconnect_2:addVector_1_avalon_rd2_read
	wire         addvector_1_avalon_rd2_readdatavalid;                         // mm_interconnect_2:addVector_1_avalon_rd2_readdatavalid -> addVector_1:masterrd2_readdatavalid
	wire   [3:0] addvector_1_avalon_rd2_burstcount;                            // addVector_1:masterrd2_burstcount -> mm_interconnect_2:addVector_1_avalon_rd2_burstcount
	wire         addvector_0_avalon_wr_waitrequest;                            // mm_interconnect_2:addVector_0_avalon_wr_waitrequest -> addVector_0:masterwr_waitrequest
	wire  [31:0] addvector_0_avalon_wr_address;                                // addVector_0:masterwr_address -> mm_interconnect_2:addVector_0_avalon_wr_address
	wire         addvector_0_avalon_wr_write;                                  // addVector_0:masterwr_write -> mm_interconnect_2:addVector_0_avalon_wr_write
	wire  [31:0] addvector_0_avalon_wr_writedata;                              // addVector_0:masterwr_writedata -> mm_interconnect_2:addVector_0_avalon_wr_writedata
	wire         addvector_1_avalon_wr_waitrequest;                            // mm_interconnect_2:addVector_1_avalon_wr_waitrequest -> addVector_1:masterwr_waitrequest
	wire  [31:0] addvector_1_avalon_wr_address;                                // addVector_1:masterwr_address -> mm_interconnect_2:addVector_1_avalon_wr_address
	wire         addvector_1_avalon_wr_write;                                  // addVector_1:masterwr_write -> mm_interconnect_2:addVector_1_avalon_wr_write
	wire  [31:0] addvector_1_avalon_wr_writedata;                              // addVector_1:masterwr_writedata -> mm_interconnect_2:addVector_1_avalon_wr_writedata
	wire  [31:0] mm_interconnect_2_hps_0_f2h_sdram0_data_readdata;             // hps_0:f2h_sdram0_READDATA -> mm_interconnect_2:hps_0_f2h_sdram0_data_readdata
	wire         mm_interconnect_2_hps_0_f2h_sdram0_data_waitrequest;          // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_2:hps_0_f2h_sdram0_data_waitrequest
	wire  [29:0] mm_interconnect_2_hps_0_f2h_sdram0_data_address;              // mm_interconnect_2:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire         mm_interconnect_2_hps_0_f2h_sdram0_data_read;                 // mm_interconnect_2:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	wire   [3:0] mm_interconnect_2_hps_0_f2h_sdram0_data_byteenable;           // mm_interconnect_2:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire         mm_interconnect_2_hps_0_f2h_sdram0_data_readdatavalid;        // hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_2:hps_0_f2h_sdram0_data_readdatavalid
	wire         mm_interconnect_2_hps_0_f2h_sdram0_data_write;                // mm_interconnect_2:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire  [31:0] mm_interconnect_2_hps_0_f2h_sdram0_data_writedata;            // mm_interconnect_2:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire   [7:0] mm_interconnect_2_hps_0_f2h_sdram0_data_burstcount;           // mm_interconnect_2:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                 // hps_0:h2f_AWBURST -> mm_interconnect_3:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                   // hps_0:h2f_ARLEN -> mm_interconnect_3:hps_0_h2f_axi_master_arlen
	wire   [7:0] hps_0_h2f_axi_master_wstrb;                                   // hps_0:h2f_WSTRB -> mm_interconnect_3:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                                  // mm_interconnect_3:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                                     // mm_interconnect_3:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                                  // hps_0:h2f_RREADY -> mm_interconnect_3:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                   // hps_0:h2f_AWLEN -> mm_interconnect_3:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                                     // hps_0:h2f_WID -> mm_interconnect_3:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                 // hps_0:h2f_ARCACHE -> mm_interconnect_3:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                                  // hps_0:h2f_WVALID -> mm_interconnect_3:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                  // hps_0:h2f_ARADDR -> mm_interconnect_3:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                  // hps_0:h2f_ARPROT -> mm_interconnect_3:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                  // hps_0:h2f_AWPROT -> mm_interconnect_3:hps_0_h2f_axi_master_awprot
	wire  [63:0] hps_0_h2f_axi_master_wdata;                                   // hps_0:h2f_WDATA -> mm_interconnect_3:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                                 // hps_0:h2f_ARVALID -> mm_interconnect_3:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                 // hps_0:h2f_AWCACHE -> mm_interconnect_3:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                                    // hps_0:h2f_ARID -> mm_interconnect_3:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                  // hps_0:h2f_ARLOCK -> mm_interconnect_3:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                  // hps_0:h2f_AWLOCK -> mm_interconnect_3:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                  // hps_0:h2f_AWADDR -> mm_interconnect_3:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                   // mm_interconnect_3:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                                 // mm_interconnect_3:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [63:0] hps_0_h2f_axi_master_rdata;                                   // mm_interconnect_3:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                                 // mm_interconnect_3:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                 // hps_0:h2f_ARBURST -> mm_interconnect_3:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                  // hps_0:h2f_ARSIZE -> mm_interconnect_3:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                                  // hps_0:h2f_BREADY -> mm_interconnect_3:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                                   // mm_interconnect_3:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                                   // hps_0:h2f_WLAST -> mm_interconnect_3:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                   // mm_interconnect_3:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                                    // hps_0:h2f_AWID -> mm_interconnect_3:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                                     // mm_interconnect_3:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                                  // mm_interconnect_3:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                  // hps_0:h2f_AWSIZE -> mm_interconnect_3:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                                 // hps_0:h2f_AWVALID -> mm_interconnect_3:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                                  // mm_interconnect_3:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_3_onchip_memory2_0_s1_chipselect;             // mm_interconnect_3:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_3_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_3:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_3_onchip_memory2_0_s1_address;                // mm_interconnect_3:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_3_onchip_memory2_0_s1_byteenable;             // mm_interconnect_3:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_3_onchip_memory2_0_s1_write;                  // mm_interconnect_3:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_3_onchip_memory2_0_s1_writedata;              // mm_interconnect_3:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_3_onchip_memory2_0_s1_clken;                  // mm_interconnect_3:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                              // hps_0:h2f_lw_AWBURST -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                // hps_0:h2f_lw_ARLEN -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                // hps_0:h2f_lw_WSTRB -> mm_interconnect_4:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                               // mm_interconnect_4:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                  // mm_interconnect_4:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                               // hps_0:h2f_lw_RREADY -> mm_interconnect_4:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                // hps_0:h2f_lw_AWLEN -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                  // hps_0:h2f_lw_WID -> mm_interconnect_4:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                              // hps_0:h2f_lw_ARCACHE -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                               // hps_0:h2f_lw_WVALID -> mm_interconnect_4:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                               // hps_0:h2f_lw_ARADDR -> mm_interconnect_4:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                               // hps_0:h2f_lw_ARPROT -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                               // hps_0:h2f_lw_AWPROT -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                // hps_0:h2f_lw_WDATA -> mm_interconnect_4:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                              // hps_0:h2f_lw_ARVALID -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                              // hps_0:h2f_lw_AWCACHE -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                 // hps_0:h2f_lw_ARID -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                               // hps_0:h2f_lw_ARLOCK -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                               // hps_0:h2f_lw_AWLOCK -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                               // hps_0:h2f_lw_AWADDR -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                // mm_interconnect_4:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                              // mm_interconnect_4:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                // mm_interconnect_4:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                              // mm_interconnect_4:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                              // hps_0:h2f_lw_ARBURST -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                               // hps_0:h2f_lw_ARSIZE -> mm_interconnect_4:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                               // hps_0:h2f_lw_BREADY -> mm_interconnect_4:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                // mm_interconnect_4:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                // hps_0:h2f_lw_WLAST -> mm_interconnect_4:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                // mm_interconnect_4:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                 // hps_0:h2f_lw_AWID -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                  // mm_interconnect_4:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                               // mm_interconnect_4:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                               // hps_0:h2f_lw_AWSIZE -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                              // hps_0:h2f_lw_AWVALID -> mm_interconnect_4:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                               // mm_interconnect_4:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_4_led_s1_chipselect;                          // mm_interconnect_4:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_4_led_s1_readdata;                            // led:readdata -> mm_interconnect_4:led_s1_readdata
	wire   [1:0] mm_interconnect_4_led_s1_address;                             // mm_interconnect_4:led_s1_address -> led:address
	wire         mm_interconnect_4_led_s1_write;                               // mm_interconnect_4:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_4_led_s1_writedata;                           // mm_interconnect_4:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_4_sw_s1_readdata;                             // sw:readdata -> mm_interconnect_4:sw_s1_readdata
	wire   [1:0] mm_interconnect_4_sw_s1_address;                              // mm_interconnect_4:sw_s1_address -> sw:address
	wire         mm_interconnect_4_bridge_stsrcmmmaster_0_slave_chipselect;    // mm_interconnect_4:bridge_stSrcMmMaster_0_slave_chipselect -> bridge_stSrcMmMaster_0:slave_chipselect
	wire  [31:0] mm_interconnect_4_bridge_stsrcmmmaster_0_slave_readdata;      // bridge_stSrcMmMaster_0:slave_readdata -> mm_interconnect_4:bridge_stSrcMmMaster_0_slave_readdata
	wire         mm_interconnect_4_bridge_stsrcmmmaster_0_slave_waitrequest;   // bridge_stSrcMmMaster_0:slave_waitrequest -> mm_interconnect_4:bridge_stSrcMmMaster_0_slave_waitrequest
	wire   [0:0] mm_interconnect_4_bridge_stsrcmmmaster_0_slave_address;       // mm_interconnect_4:bridge_stSrcMmMaster_0_slave_address -> bridge_stSrcMmMaster_0:slave_address
	wire         mm_interconnect_4_bridge_stsrcmmmaster_0_slave_read;          // mm_interconnect_4:bridge_stSrcMmMaster_0_slave_read -> bridge_stSrcMmMaster_0:slave_read
	wire         mm_interconnect_4_bridge_stsrcmmmaster_0_slave_readdatavalid; // bridge_stSrcMmMaster_0:slave_readdatavalid -> mm_interconnect_4:bridge_stSrcMmMaster_0_slave_readdatavalid
	wire         mm_interconnect_4_bridge_stsrcmmmaster_0_slave_write;         // mm_interconnect_4:bridge_stSrcMmMaster_0_slave_write -> bridge_stSrcMmMaster_0:slave_write
	wire  [31:0] mm_interconnect_4_bridge_stsrcmmmaster_0_slave_writedata;     // mm_interconnect_4:bridge_stSrcMmMaster_0_slave_writedata -> bridge_stSrcMmMaster_0:slave_writedata
	wire         mm_interconnect_4_lwir_ul0304_0_slave_chipselect;             // mm_interconnect_4:lwir_ul0304_0_slave_chipselect -> lwir_ul0304_0:slave_chipselect
	wire  [31:0] mm_interconnect_4_lwir_ul0304_0_slave_readdata;               // lwir_ul0304_0:slave_readdata -> mm_interconnect_4:lwir_ul0304_0_slave_readdata
	wire         mm_interconnect_4_lwir_ul0304_0_slave_waitrequest;            // lwir_ul0304_0:slave_waitrequest -> mm_interconnect_4:lwir_ul0304_0_slave_waitrequest
	wire   [0:0] mm_interconnect_4_lwir_ul0304_0_slave_address;                // mm_interconnect_4:lwir_ul0304_0_slave_address -> lwir_ul0304_0:slave_address
	wire         mm_interconnect_4_lwir_ul0304_0_slave_read;                   // mm_interconnect_4:lwir_ul0304_0_slave_read -> lwir_ul0304_0:slave_read
	wire   [3:0] mm_interconnect_4_lwir_ul0304_0_slave_byteenable;             // mm_interconnect_4:lwir_ul0304_0_slave_byteenable -> lwir_ul0304_0:slave_byteenable
	wire         mm_interconnect_4_lwir_ul0304_0_slave_readdatavalid;          // lwir_ul0304_0:slave_readdatavalid -> mm_interconnect_4:lwir_ul0304_0_slave_readdatavalid
	wire         mm_interconnect_4_lwir_ul0304_0_slave_write;                  // mm_interconnect_4:lwir_ul0304_0_slave_write -> lwir_ul0304_0:slave_write
	wire  [31:0] mm_interconnect_4_lwir_ul0304_0_slave_writedata;              // mm_interconnect_4:lwir_ul0304_0_slave_writedata -> lwir_ul0304_0:slave_writedata
	wire         mm_interconnect_4_swir_v400_0_slave_chipselect;               // mm_interconnect_4:swir_v400_0_slave_chipselect -> swir_v400_0:slave_chipselect
	wire  [31:0] mm_interconnect_4_swir_v400_0_slave_readdata;                 // swir_v400_0:slave_readdata -> mm_interconnect_4:swir_v400_0_slave_readdata
	wire         mm_interconnect_4_swir_v400_0_slave_waitrequest;              // swir_v400_0:slave_waitrequest -> mm_interconnect_4:swir_v400_0_slave_waitrequest
	wire   [0:0] mm_interconnect_4_swir_v400_0_slave_address;                  // mm_interconnect_4:swir_v400_0_slave_address -> swir_v400_0:slave_address
	wire         mm_interconnect_4_swir_v400_0_slave_read;                     // mm_interconnect_4:swir_v400_0_slave_read -> swir_v400_0:slave_read
	wire   [3:0] mm_interconnect_4_swir_v400_0_slave_byteenable;               // mm_interconnect_4:swir_v400_0_slave_byteenable -> swir_v400_0:slave_byteenable
	wire         mm_interconnect_4_swir_v400_0_slave_readdatavalid;            // swir_v400_0:slave_readdatavalid -> mm_interconnect_4:swir_v400_0_slave_readdatavalid
	wire         mm_interconnect_4_swir_v400_0_slave_write;                    // mm_interconnect_4:swir_v400_0_slave_write -> swir_v400_0:slave_write
	wire  [31:0] mm_interconnect_4_swir_v400_0_slave_writedata;                // mm_interconnect_4:swir_v400_0_slave_writedata -> swir_v400_0:slave_writedata
	wire         mm_interconnect_4_bridge_stsrcmmmaster_1_slave_chipselect;    // mm_interconnect_4:bridge_stSrcMmMaster_1_slave_chipselect -> bridge_stSrcMmMaster_1:slave_chipselect
	wire  [31:0] mm_interconnect_4_bridge_stsrcmmmaster_1_slave_readdata;      // bridge_stSrcMmMaster_1:slave_readdata -> mm_interconnect_4:bridge_stSrcMmMaster_1_slave_readdata
	wire         mm_interconnect_4_bridge_stsrcmmmaster_1_slave_waitrequest;   // bridge_stSrcMmMaster_1:slave_waitrequest -> mm_interconnect_4:bridge_stSrcMmMaster_1_slave_waitrequest
	wire   [0:0] mm_interconnect_4_bridge_stsrcmmmaster_1_slave_address;       // mm_interconnect_4:bridge_stSrcMmMaster_1_slave_address -> bridge_stSrcMmMaster_1:slave_address
	wire         mm_interconnect_4_bridge_stsrcmmmaster_1_slave_read;          // mm_interconnect_4:bridge_stSrcMmMaster_1_slave_read -> bridge_stSrcMmMaster_1:slave_read
	wire         mm_interconnect_4_bridge_stsrcmmmaster_1_slave_readdatavalid; // bridge_stSrcMmMaster_1:slave_readdatavalid -> mm_interconnect_4:bridge_stSrcMmMaster_1_slave_readdatavalid
	wire         mm_interconnect_4_bridge_stsrcmmmaster_1_slave_write;         // mm_interconnect_4:bridge_stSrcMmMaster_1_slave_write -> bridge_stSrcMmMaster_1:slave_write
	wire  [31:0] mm_interconnect_4_bridge_stsrcmmmaster_1_slave_writedata;     // mm_interconnect_4:bridge_stSrcMmMaster_1_slave_writedata -> bridge_stSrcMmMaster_1:slave_writedata
	wire         mm_interconnect_4_addvector_0_slave_1_chipselect;             // mm_interconnect_4:addVector_0_slave_1_chipselect -> addVector_0:slave_chipselect
	wire  [31:0] mm_interconnect_4_addvector_0_slave_1_readdata;               // addVector_0:slave_readdata -> mm_interconnect_4:addVector_0_slave_1_readdata
	wire         mm_interconnect_4_addvector_0_slave_1_waitrequest;            // addVector_0:slave_waitrequest -> mm_interconnect_4:addVector_0_slave_1_waitrequest
	wire   [2:0] mm_interconnect_4_addvector_0_slave_1_address;                // mm_interconnect_4:addVector_0_slave_1_address -> addVector_0:slave_address
	wire         mm_interconnect_4_addvector_0_slave_1_read;                   // mm_interconnect_4:addVector_0_slave_1_read -> addVector_0:slave_read
	wire   [3:0] mm_interconnect_4_addvector_0_slave_1_byteenable;             // mm_interconnect_4:addVector_0_slave_1_byteenable -> addVector_0:slave_byteenable
	wire         mm_interconnect_4_addvector_0_slave_1_readdatavalid;          // addVector_0:slave_readdatavalid -> mm_interconnect_4:addVector_0_slave_1_readdatavalid
	wire         mm_interconnect_4_addvector_0_slave_1_write;                  // mm_interconnect_4:addVector_0_slave_1_write -> addVector_0:slave_write
	wire  [31:0] mm_interconnect_4_addvector_0_slave_1_writedata;              // mm_interconnect_4:addVector_0_slave_1_writedata -> addVector_0:slave_writedata
	wire         mm_interconnect_4_addvector_1_slave_1_chipselect;             // mm_interconnect_4:addVector_1_slave_1_chipselect -> addVector_1:slave_chipselect
	wire  [31:0] mm_interconnect_4_addvector_1_slave_1_readdata;               // addVector_1:slave_readdata -> mm_interconnect_4:addVector_1_slave_1_readdata
	wire         mm_interconnect_4_addvector_1_slave_1_waitrequest;            // addVector_1:slave_waitrequest -> mm_interconnect_4:addVector_1_slave_1_waitrequest
	wire   [2:0] mm_interconnect_4_addvector_1_slave_1_address;                // mm_interconnect_4:addVector_1_slave_1_address -> addVector_1:slave_address
	wire         mm_interconnect_4_addvector_1_slave_1_read;                   // mm_interconnect_4:addVector_1_slave_1_read -> addVector_1:slave_read
	wire   [3:0] mm_interconnect_4_addvector_1_slave_1_byteenable;             // mm_interconnect_4:addVector_1_slave_1_byteenable -> addVector_1:slave_byteenable
	wire         mm_interconnect_4_addvector_1_slave_1_readdatavalid;          // addVector_1:slave_readdatavalid -> mm_interconnect_4:addVector_1_slave_1_readdatavalid
	wire         mm_interconnect_4_addvector_1_slave_1_write;                  // mm_interconnect_4:addVector_1_slave_1_write -> addVector_1:slave_write
	wire  [31:0] mm_interconnect_4_addvector_1_slave_1_writedata;              // mm_interconnect_4:addVector_1_slave_1_writedata -> addVector_1:slave_writedata
	wire         lwir_ul0304_0_st_valid;                                       // lwir_ul0304_0:st_data_valid -> avalon_st_adapter:in_0_valid
	wire   [7:0] lwir_ul0304_0_st_data;                                        // lwir_ul0304_0:st_data_out -> avalon_st_adapter:in_0_data
	wire         lwir_ul0304_0_st_startofpacket;                               // lwir_ul0304_0:st_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         lwir_ul0304_0_st_endofpacket;                                 // lwir_ul0304_0:st_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                // avalon_st_adapter:out_0_valid -> bridge_stSrcMmMaster_0:st_datavalid
	wire   [7:0] avalon_st_adapter_out_0_data;                                 // avalon_st_adapter:out_0_data -> bridge_stSrcMmMaster_0:st_datain
	wire         avalon_st_adapter_out_0_ready;                                // bridge_stSrcMmMaster_0:st_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                        // avalon_st_adapter:out_0_startofpacket -> bridge_stSrcMmMaster_0:st_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                          // avalon_st_adapter:out_0_endofpacket -> bridge_stSrcMmMaster_0:st_endofpacket
	wire         swir_v400_0_st_valid;                                         // swir_v400_0:st_data_valid -> avalon_st_adapter_001:in_0_valid
	wire   [7:0] swir_v400_0_st_data;                                          // swir_v400_0:st_data_out -> avalon_st_adapter_001:in_0_data
	wire         swir_v400_0_st_startofpacket;                                 // swir_v400_0:st_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire         swir_v400_0_st_endofpacket;                                   // swir_v400_0:st_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;                            // avalon_st_adapter_001:out_0_valid -> bridge_stSrcMmMaster_1:st_datavalid
	wire   [7:0] avalon_st_adapter_001_out_0_data;                             // avalon_st_adapter_001:out_0_data -> bridge_stSrcMmMaster_1:st_datain
	wire         avalon_st_adapter_001_out_0_ready;                            // bridge_stSrcMmMaster_1:st_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;                    // avalon_st_adapter_001:out_0_startofpacket -> bridge_stSrcMmMaster_1:st_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                      // avalon_st_adapter_001:out_0_endofpacket -> bridge_stSrcMmMaster_1:st_endofpacket
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [addVector_0:rst_n, addVector_1:rst_n, led:reset_n, mm_interconnect_0:bridge_stSrcMmMaster_1_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:bridge_stSrcMmMaster_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:addVector_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_3:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_4:led_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, sw:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, bridge_stSrcMmMaster_0:rst_n, lwir_ul0304_0:rst_n, mm_interconnect_4:lwir_ul0304_0_reset_sink_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [avalon_st_adapter_001:in_rst_0_reset, bridge_stSrcMmMaster_1:rst_n, mm_interconnect_4:swir_v400_0_reset_sink_reset_bridge_in_reset_reset, swir_v400_0:rst_n]
	wire         rst_controller_003_reset_out_reset;                           // rst_controller_003:reset_out -> [mm_interconnect_0:hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_f2h_sdram3_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_4:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire         hps_0_h2f_reset_reset;                                        // hps_0:h2f_rst_n -> rst_controller_003:reset_in0

	addVector_avalon #(
		.NBITS_ADDR    (32),
		.NBITS_PACKETS (32),
		.FIFO_SIZE     (256),
		.NBITS_DATA    (32),
		.NBITS_BURST   (4),
		.NBITS_BYTEEN  (4),
		.BURST         (8),
		.ADDR_READ1    (32'b00111000000000000000000000000000),
		.ADDR_READ2    (32'b00111000000100000000000000000000),
		.ADDR_WRITE    (32'b00111000110000000000000000000000)
	) addvector_0 (
		.clk                     (clk_clk),                                             //            clock.clk
		.rst_n                   (~rst_controller_reset_out_reset),                     //       reset_sink.reset_n
		.slave_chipselect        (mm_interconnect_4_addvector_0_slave_1_chipselect),    //          slave_1.chipselect
		.slave_read              (mm_interconnect_4_addvector_0_slave_1_read),          //                 .read
		.slave_write             (mm_interconnect_4_addvector_0_slave_1_write),         //                 .write
		.slave_address           (mm_interconnect_4_addvector_0_slave_1_address),       //                 .address
		.slave_writedata         (mm_interconnect_4_addvector_0_slave_1_writedata),     //                 .writedata
		.slave_waitrequest       (mm_interconnect_4_addvector_0_slave_1_waitrequest),   //                 .waitrequest
		.slave_readdatavalid     (mm_interconnect_4_addvector_0_slave_1_readdatavalid), //                 .readdatavalid
		.slave_readdata          (mm_interconnect_4_addvector_0_slave_1_readdata),      //                 .readdata
		.slave_byteenable        (mm_interconnect_4_addvector_0_slave_1_byteenable),    //                 .byteenable
		.masterwr_address        (addvector_0_avalon_wr_address),                       //        avalon_wr.address
		.masterwr_waitrequest    (addvector_0_avalon_wr_waitrequest),                   //                 .waitrequest
		.masterwr_write          (addvector_0_avalon_wr_write),                         //                 .write
		.masterwr_writedata      (addvector_0_avalon_wr_writedata),                     //                 .writedata
		.masterrd2_address       (addvector_0_avalon_rd2_address),                      //       avalon_rd2.address
		.masterrd2_read          (addvector_0_avalon_rd2_read),                         //                 .read
		.masterrd2_readdata      (addvector_0_avalon_rd2_readdata),                     //                 .readdata
		.masterrd2_readdatavalid (addvector_0_avalon_rd2_readdatavalid),                //                 .readdatavalid
		.masterrd2_waitrequest   (addvector_0_avalon_rd2_waitrequest),                  //                 .waitrequest
		.masterrd2_burstcount    (addvector_0_avalon_rd2_burstcount),                   //                 .burstcount
		.masterrd1_address       (addvector_0_avalon_rd1_1_1_1_address),                // avalon_rd1_1_1_1.address
		.masterrd1_read          (addvector_0_avalon_rd1_1_1_1_read),                   //                 .read
		.masterrd1_readdata      (addvector_0_avalon_rd1_1_1_1_readdata),               //                 .readdata
		.masterrd1_readdatavalid (addvector_0_avalon_rd1_1_1_1_readdatavalid),          //                 .readdatavalid
		.masterrd1_waitrequest   (addvector_0_avalon_rd1_1_1_1_waitrequest),            //                 .waitrequest
		.masterrd1_burstcount    (addvector_0_avalon_rd1_1_1_1_burstcount)              //                 .burstcount
	);

	addVector_avalon #(
		.NBITS_ADDR    (32),
		.NBITS_PACKETS (32),
		.FIFO_SIZE     (256),
		.NBITS_DATA    (32),
		.NBITS_BURST   (4),
		.NBITS_BYTEEN  (4),
		.BURST         (8),
		.ADDR_READ1    (32'b00111000001000000000000000000000),
		.ADDR_READ2    (32'b00111000001100000000000000000000),
		.ADDR_WRITE    (32'b00111000010000000000000000000000)
	) addvector_1 (
		.clk                     (clk_clk),                                             //            clock.clk
		.rst_n                   (~rst_controller_reset_out_reset),                     //       reset_sink.reset_n
		.slave_chipselect        (mm_interconnect_4_addvector_1_slave_1_chipselect),    //          slave_1.chipselect
		.slave_read              (mm_interconnect_4_addvector_1_slave_1_read),          //                 .read
		.slave_write             (mm_interconnect_4_addvector_1_slave_1_write),         //                 .write
		.slave_address           (mm_interconnect_4_addvector_1_slave_1_address),       //                 .address
		.slave_writedata         (mm_interconnect_4_addvector_1_slave_1_writedata),     //                 .writedata
		.slave_waitrequest       (mm_interconnect_4_addvector_1_slave_1_waitrequest),   //                 .waitrequest
		.slave_readdatavalid     (mm_interconnect_4_addvector_1_slave_1_readdatavalid), //                 .readdatavalid
		.slave_readdata          (mm_interconnect_4_addvector_1_slave_1_readdata),      //                 .readdata
		.slave_byteenable        (mm_interconnect_4_addvector_1_slave_1_byteenable),    //                 .byteenable
		.masterwr_address        (addvector_1_avalon_wr_address),                       //        avalon_wr.address
		.masterwr_waitrequest    (addvector_1_avalon_wr_waitrequest),                   //                 .waitrequest
		.masterwr_write          (addvector_1_avalon_wr_write),                         //                 .write
		.masterwr_writedata      (addvector_1_avalon_wr_writedata),                     //                 .writedata
		.masterrd2_address       (addvector_1_avalon_rd2_address),                      //       avalon_rd2.address
		.masterrd2_read          (addvector_1_avalon_rd2_read),                         //                 .read
		.masterrd2_readdata      (addvector_1_avalon_rd2_readdata),                     //                 .readdata
		.masterrd2_readdatavalid (addvector_1_avalon_rd2_readdatavalid),                //                 .readdatavalid
		.masterrd2_waitrequest   (addvector_1_avalon_rd2_waitrequest),                  //                 .waitrequest
		.masterrd2_burstcount    (addvector_1_avalon_rd2_burstcount),                   //                 .burstcount
		.masterrd1_address       (addvector_1_avalon_rd1_1_1_1_address),                // avalon_rd1_1_1_1.address
		.masterrd1_read          (addvector_1_avalon_rd1_1_1_1_read),                   //                 .read
		.masterrd1_readdata      (addvector_1_avalon_rd1_1_1_1_readdata),               //                 .readdata
		.masterrd1_readdatavalid (addvector_1_avalon_rd1_1_1_1_readdatavalid),          //                 .readdatavalid
		.masterrd1_waitrequest   (addvector_1_avalon_rd1_1_1_1_waitrequest),            //                 .waitrequest
		.masterrd1_burstcount    (addvector_1_avalon_rd1_1_1_1_burstcount)              //                 .burstcount
	);

	bridge_stSrc_mmMaster #(
		.NBITS_ADDR    (32),
		.NBITS_DATA    (8),
		.NBITS_BURST   (4),
		.NBITS_BYTEEN  (4),
		.BURST         (1),
		.ADDR_BASE_BUF (32'b00111000000000000000000000000000)
	) bridge_stsrcmmmaster_0 (
		.clk                 (pll_0_outclk1_clk),                                            //                 clock.clk
		.master_waitrequest  (bridge_stsrcmmmaster_0_avalon_master_waitrequest),             //         avalon_master.waitrequest
		.master_address      (bridge_stsrcmmmaster_0_avalon_master_address),                 //                      .address
		.master_write        (bridge_stsrcmmmaster_0_avalon_master_write),                   //                      .write
		.master_writedata    (bridge_stsrcmmmaster_0_avalon_master_writedata),               //                      .writedata
		.master_burstcount   (bridge_stsrcmmmaster_0_avalon_master_burstcount),              //                      .burstcount
		.st_datain           (avalon_st_adapter_out_0_data),                                 // avalon_streaming_sink.data
		.st_datavalid        (avalon_st_adapter_out_0_valid),                                //                      .valid
		.st_endofpacket      (avalon_st_adapter_out_0_endofpacket),                          //                      .endofpacket
		.st_ready            (avalon_st_adapter_out_0_ready),                                //                      .ready
		.st_startofpacket    (avalon_st_adapter_out_0_startofpacket),                        //                      .startofpacket
		.rst_n               (~rst_controller_001_reset_out_reset),                          //            reset_sink.reset_n
		.clk_mem             (clk_clk),                                                      //             clock_mem.clk
		.slave_chipselect    (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_chipselect),    //                 slave.chipselect
		.slave_read          (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_read),          //                      .read
		.slave_write         (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_write),         //                      .write
		.slave_address       (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_address),       //                      .address
		.slave_writedata     (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_writedata),     //                      .writedata
		.slave_waitrequest   (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_waitrequest),   //                      .waitrequest
		.slave_readdatavalid (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_readdatavalid), //                      .readdatavalid
		.slave_readdata      (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_readdata)       //                      .readdata
	);

	bridge_stSrc_mmMaster #(
		.NBITS_ADDR    (32),
		.NBITS_DATA    (8),
		.NBITS_BURST   (4),
		.NBITS_BYTEEN  (4),
		.BURST         (1),
		.ADDR_BASE_BUF (32'b00111000001000000000000000000000)
	) bridge_stsrcmmmaster_1 (
		.clk                 (pll_0_outclk0_clk),                                            //                 clock.clk
		.master_waitrequest  (bridge_stsrcmmmaster_1_avalon_master_waitrequest),             //         avalon_master.waitrequest
		.master_address      (bridge_stsrcmmmaster_1_avalon_master_address),                 //                      .address
		.master_write        (bridge_stsrcmmmaster_1_avalon_master_write),                   //                      .write
		.master_writedata    (bridge_stsrcmmmaster_1_avalon_master_writedata),               //                      .writedata
		.master_burstcount   (bridge_stsrcmmmaster_1_avalon_master_burstcount),              //                      .burstcount
		.st_datain           (avalon_st_adapter_001_out_0_data),                             // avalon_streaming_sink.data
		.st_datavalid        (avalon_st_adapter_001_out_0_valid),                            //                      .valid
		.st_endofpacket      (avalon_st_adapter_001_out_0_endofpacket),                      //                      .endofpacket
		.st_ready            (avalon_st_adapter_001_out_0_ready),                            //                      .ready
		.st_startofpacket    (avalon_st_adapter_001_out_0_startofpacket),                    //                      .startofpacket
		.rst_n               (~rst_controller_002_reset_out_reset),                          //            reset_sink.reset_n
		.clk_mem             (clk_clk),                                                      //             clock_mem.clk
		.slave_chipselect    (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_chipselect),    //                 slave.chipselect
		.slave_read          (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_read),          //                      .read
		.slave_write         (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_write),         //                      .write
		.slave_address       (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_address),       //                      .address
		.slave_writedata     (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_writedata),     //                      .writedata
		.slave_waitrequest   (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_waitrequest),   //                      .waitrequest
		.slave_readdatavalid (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_readdatavalid), //                      .readdatavalid
		.slave_readdata      (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_readdata)       //                      .readdata
	);

	cycloneV_soc_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                          //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                         //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                         //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                       //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                        //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                       //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                      //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                      //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                       //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                    //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                         //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                        //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                      //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                        //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                         //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                      //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                       //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                         //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                         //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                         //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                         //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                         //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                         //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                          //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                       //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                       //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                       //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                         //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                         //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                         //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                           //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                            //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                            //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                           //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                            //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                            //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                            //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                            //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                            //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                            //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                            //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                            //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                            //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                            //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                           //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                           //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                           //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                           //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                           //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                           //                  .hps_io_uart0_inst_TX
		.h2f_rst_n                (hps_0_h2f_reset_reset),                                 //         h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                                               //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_2_hps_0_f2h_sdram0_data_address),       //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_2_hps_0_f2h_sdram0_data_burstcount),    //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_2_hps_0_f2h_sdram0_data_waitrequest),   //                  .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_2_hps_0_f2h_sdram0_data_readdata),      //                  .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_2_hps_0_f2h_sdram0_data_readdatavalid), //                  .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_2_hps_0_f2h_sdram0_data_read),          //                  .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_2_hps_0_f2h_sdram0_data_writedata),     //                  .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_2_hps_0_f2h_sdram0_data_byteenable),    //                  .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_2_hps_0_f2h_sdram0_data_write),         //                  .write
		.f2h_sdram1_clk           (clk_clk),                                               //  f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS       (mm_interconnect_0_hps_0_f2h_sdram1_data_address),       //   f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT    (mm_interconnect_0_hps_0_f2h_sdram1_data_burstcount),    //                  .burstcount
		.f2h_sdram1_WAITREQUEST   (mm_interconnect_0_hps_0_f2h_sdram1_data_waitrequest),   //                  .waitrequest
		.f2h_sdram1_WRITEDATA     (mm_interconnect_0_hps_0_f2h_sdram1_data_writedata),     //                  .writedata
		.f2h_sdram1_BYTEENABLE    (mm_interconnect_0_hps_0_f2h_sdram1_data_byteenable),    //                  .byteenable
		.f2h_sdram1_WRITE         (mm_interconnect_0_hps_0_f2h_sdram1_data_write),         //                  .write
		.f2h_sdram2_clk           (clk_clk),                                               //  f2h_sdram2_clock.clk
		.f2h_sdram2_ADDRESS       (),                                                      //   f2h_sdram2_data.address
		.f2h_sdram2_BURSTCOUNT    (),                                                      //                  .burstcount
		.f2h_sdram2_WAITREQUEST   (),                                                      //                  .waitrequest
		.f2h_sdram2_READDATA      (),                                                      //                  .readdata
		.f2h_sdram2_READDATAVALID (),                                                      //                  .readdatavalid
		.f2h_sdram2_READ          (),                                                      //                  .read
		.f2h_sdram2_WRITEDATA     (),                                                      //                  .writedata
		.f2h_sdram2_BYTEENABLE    (),                                                      //                  .byteenable
		.f2h_sdram2_WRITE         (),                                                      //                  .write
		.f2h_sdram3_clk           (clk_clk),                                               //  f2h_sdram3_clock.clk
		.f2h_sdram3_ADDRESS       (mm_interconnect_1_hps_0_f2h_sdram3_data_address),       //   f2h_sdram3_data.address
		.f2h_sdram3_BURSTCOUNT    (mm_interconnect_1_hps_0_f2h_sdram3_data_burstcount),    //                  .burstcount
		.f2h_sdram3_WAITREQUEST   (mm_interconnect_1_hps_0_f2h_sdram3_data_waitrequest),   //                  .waitrequest
		.f2h_sdram3_WRITEDATA     (mm_interconnect_1_hps_0_f2h_sdram3_data_writedata),     //                  .writedata
		.f2h_sdram3_BYTEENABLE    (mm_interconnect_1_hps_0_f2h_sdram3_data_byteenable),    //                  .byteenable
		.f2h_sdram3_WRITE         (mm_interconnect_1_hps_0_f2h_sdram3_data_write),         //                  .write
		.h2f_axi_clk              (clk_clk),                                               //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                             //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                           //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                            //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                           //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                          //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                           //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                          //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                           //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                          //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                          //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                              //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                            //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                            //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                            //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                           //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                           //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                              //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                            //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                           //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                           //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                             //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                           //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                            //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                           //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                          //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                           //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                          //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                           //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                          //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                          //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                              //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                            //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                            //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                            //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                           //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                           //                  .rready
		.f2h_axi_clk              (clk_clk),                                               //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                                      //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                      //                  .awaddr
		.f2h_AWLEN                (),                                                      //                  .awlen
		.f2h_AWSIZE               (),                                                      //                  .awsize
		.f2h_AWBURST              (),                                                      //                  .awburst
		.f2h_AWLOCK               (),                                                      //                  .awlock
		.f2h_AWCACHE              (),                                                      //                  .awcache
		.f2h_AWPROT               (),                                                      //                  .awprot
		.f2h_AWVALID              (),                                                      //                  .awvalid
		.f2h_AWREADY              (),                                                      //                  .awready
		.f2h_AWUSER               (),                                                      //                  .awuser
		.f2h_WID                  (),                                                      //                  .wid
		.f2h_WDATA                (),                                                      //                  .wdata
		.f2h_WSTRB                (),                                                      //                  .wstrb
		.f2h_WLAST                (),                                                      //                  .wlast
		.f2h_WVALID               (),                                                      //                  .wvalid
		.f2h_WREADY               (),                                                      //                  .wready
		.f2h_BID                  (),                                                      //                  .bid
		.f2h_BRESP                (),                                                      //                  .bresp
		.f2h_BVALID               (),                                                      //                  .bvalid
		.f2h_BREADY               (),                                                      //                  .bready
		.f2h_ARID                 (),                                                      //                  .arid
		.f2h_ARADDR               (),                                                      //                  .araddr
		.f2h_ARLEN                (),                                                      //                  .arlen
		.f2h_ARSIZE               (),                                                      //                  .arsize
		.f2h_ARBURST              (),                                                      //                  .arburst
		.f2h_ARLOCK               (),                                                      //                  .arlock
		.f2h_ARCACHE              (),                                                      //                  .arcache
		.f2h_ARPROT               (),                                                      //                  .arprot
		.f2h_ARVALID              (),                                                      //                  .arvalid
		.f2h_ARREADY              (),                                                      //                  .arready
		.f2h_ARUSER               (),                                                      //                  .aruser
		.f2h_RID                  (),                                                      //                  .rid
		.f2h_RDATA                (),                                                      //                  .rdata
		.f2h_RRESP                (),                                                      //                  .rresp
		.f2h_RLAST                (),                                                      //                  .rlast
		.f2h_RVALID               (),                                                      //                  .rvalid
		.f2h_RREADY               (),                                                      //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                                               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                        //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                         //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                        //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                       //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                        //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                       //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                        //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                       //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                       //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                           //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                         //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                         //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                         //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                        //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                        //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                           //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                         //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                        //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                        //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                          //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                        //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                         //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                        //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                       //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                        //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                       //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                        //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                       //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                       //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                           //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                         //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                         //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                         //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                        //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)                         //                  .rready
	);

	cycloneV_soc_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_4_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_4_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_4_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_4_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_4_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	lwir_ul0304_avalon #(
		.NUM_COLS  (320),
		.NUM_ROWS  (256),
		.NBITS_PXL (8)
	) lwir_ul0304_0 (
		.slave_chipselect    (mm_interconnect_4_lwir_ul0304_0_slave_chipselect),    //       slave.chipselect
		.slave_read          (mm_interconnect_4_lwir_ul0304_0_slave_read),          //            .read
		.slave_write         (mm_interconnect_4_lwir_ul0304_0_slave_write),         //            .write
		.slave_address       (mm_interconnect_4_lwir_ul0304_0_slave_address),       //            .address
		.slave_byteenable    (mm_interconnect_4_lwir_ul0304_0_slave_byteenable),    //            .byteenable
		.slave_writedata     (mm_interconnect_4_lwir_ul0304_0_slave_writedata),     //            .writedata
		.slave_waitrequest   (mm_interconnect_4_lwir_ul0304_0_slave_waitrequest),   //            .waitrequest
		.slave_readdatavalid (mm_interconnect_4_lwir_ul0304_0_slave_readdatavalid), //            .readdatavalid
		.slave_readdata      (mm_interconnect_4_lwir_ul0304_0_slave_readdata),      //            .readdata
		.st_endofpacket      (lwir_ul0304_0_st_endofpacket),                        //          st.endofpacket
		.st_data_out         (lwir_ul0304_0_st_data),                               //            .data
		.st_data_valid       (lwir_ul0304_0_st_valid),                              //            .valid
		.st_startofpacket    (lwir_ul0304_0_st_startofpacket),                      //            .startofpacket
		.sensor_clk_in       (pll_0_outclk1_clk),                                   //  clock_sink.clk
		.rst_n               (~rst_controller_001_reset_out_reset),                 //  reset_sink.reset_n
		.lwir_dataIn         (lwir_ul0304_datain),                                  // conduit_end.datain
		.lwir_syt            (lwir_ul0304_syt),                                     //            .syt
		.lwir_syl            (lwir_ul0304_syl),                                     //            .syl
		.lwir_syp            (lwir_ul0304_syp)                                      //            .syp
	);

	cycloneV_soc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_3_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_3_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_3_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_3_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_3_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_3_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_3_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	cycloneV_soc_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.locked   ()                   //  locked.export
	);

	cycloneV_soc_sw sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_4_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_4_sw_s1_readdata), //                    .readdata
		.in_port  (sw_external_connection_export)     // external_connection.export
	);

	swir_controller_avalon swir_v400_0 (
		.slave_chipselect    (mm_interconnect_4_swir_v400_0_slave_chipselect),    //       slave.chipselect
		.slave_read          (mm_interconnect_4_swir_v400_0_slave_read),          //            .read
		.slave_write         (mm_interconnect_4_swir_v400_0_slave_write),         //            .write
		.slave_address       (mm_interconnect_4_swir_v400_0_slave_address),       //            .address
		.slave_byteenable    (mm_interconnect_4_swir_v400_0_slave_byteenable),    //            .byteenable
		.slave_writedata     (mm_interconnect_4_swir_v400_0_slave_writedata),     //            .writedata
		.slave_waitrequest   (mm_interconnect_4_swir_v400_0_slave_waitrequest),   //            .waitrequest
		.slave_readdatavalid (mm_interconnect_4_swir_v400_0_slave_readdatavalid), //            .readdatavalid
		.slave_readdata      (mm_interconnect_4_swir_v400_0_slave_readdata),      //            .readdata
		.st_endofpacket      (swir_v400_0_st_endofpacket),                        //          st.endofpacket
		.st_data_out         (swir_v400_0_st_data),                               //            .data
		.st_data_valid       (swir_v400_0_st_valid),                              //            .valid
		.st_startofpacket    (swir_v400_0_st_startofpacket),                      //            .startofpacket
		.pxl_clk_in          (pll_0_outclk0_clk),                                 //     pxl_clk.clk
		.sensor_clk_in       (pll_0_outclk1_clk),                                 //  sensor_clk.clk
		.swir_clk_out        (swir_v400_sensor_clk),                              // conduit_end.sensor_clk
		.swir_dataIn         (swir_v400_datain),                                  //            .datain
		.swir_fsync          (swir_v400_fsync),                                   //            .fsync
		.swir_lsync          (swir_v400_lsync),                                   //            .lsync
		.swir_pclk_out       (swir_v400_swir_pxl_clk_out),                        //            .swir_pxl_clk_out
		.rst_n               (~rst_controller_002_reset_out_reset)                //  reset_sink.reset_n
	);

	cycloneV_soc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                      (clk_clk),                                             //                                                    clk_0_clk.clk
		.bridge_stSrcMmMaster_1_reset_sink_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                      //      bridge_stSrcMmMaster_1_reset_sink_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                  // hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset.reset
		.bridge_stSrcMmMaster_1_avalon_master_address                       (bridge_stsrcmmmaster_1_avalon_master_address),        //                         bridge_stSrcMmMaster_1_avalon_master.address
		.bridge_stSrcMmMaster_1_avalon_master_waitrequest                   (bridge_stsrcmmmaster_1_avalon_master_waitrequest),    //                                                             .waitrequest
		.bridge_stSrcMmMaster_1_avalon_master_burstcount                    (bridge_stsrcmmmaster_1_avalon_master_burstcount),     //                                                             .burstcount
		.bridge_stSrcMmMaster_1_avalon_master_write                         (bridge_stsrcmmmaster_1_avalon_master_write),          //                                                             .write
		.bridge_stSrcMmMaster_1_avalon_master_writedata                     (bridge_stsrcmmmaster_1_avalon_master_writedata),      //                                                             .writedata
		.hps_0_f2h_sdram1_data_address                                      (mm_interconnect_0_hps_0_f2h_sdram1_data_address),     //                                        hps_0_f2h_sdram1_data.address
		.hps_0_f2h_sdram1_data_write                                        (mm_interconnect_0_hps_0_f2h_sdram1_data_write),       //                                                             .write
		.hps_0_f2h_sdram1_data_writedata                                    (mm_interconnect_0_hps_0_f2h_sdram1_data_writedata),   //                                                             .writedata
		.hps_0_f2h_sdram1_data_burstcount                                   (mm_interconnect_0_hps_0_f2h_sdram1_data_burstcount),  //                                                             .burstcount
		.hps_0_f2h_sdram1_data_byteenable                                   (mm_interconnect_0_hps_0_f2h_sdram1_data_byteenable),  //                                                             .byteenable
		.hps_0_f2h_sdram1_data_waitrequest                                  (mm_interconnect_0_hps_0_f2h_sdram1_data_waitrequest)  //                                                             .waitrequest
	);

	cycloneV_soc_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                                      (clk_clk),                                             //                                                    clk_0_clk.clk
		.bridge_stSrcMmMaster_0_reset_sink_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                      //      bridge_stSrcMmMaster_0_reset_sink_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram3_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                  // hps_0_f2h_sdram3_data_translator_reset_reset_bridge_in_reset.reset
		.bridge_stSrcMmMaster_0_avalon_master_address                       (bridge_stsrcmmmaster_0_avalon_master_address),        //                         bridge_stSrcMmMaster_0_avalon_master.address
		.bridge_stSrcMmMaster_0_avalon_master_waitrequest                   (bridge_stsrcmmmaster_0_avalon_master_waitrequest),    //                                                             .waitrequest
		.bridge_stSrcMmMaster_0_avalon_master_burstcount                    (bridge_stsrcmmmaster_0_avalon_master_burstcount),     //                                                             .burstcount
		.bridge_stSrcMmMaster_0_avalon_master_write                         (bridge_stsrcmmmaster_0_avalon_master_write),          //                                                             .write
		.bridge_stSrcMmMaster_0_avalon_master_writedata                     (bridge_stsrcmmmaster_0_avalon_master_writedata),      //                                                             .writedata
		.hps_0_f2h_sdram3_data_address                                      (mm_interconnect_1_hps_0_f2h_sdram3_data_address),     //                                        hps_0_f2h_sdram3_data.address
		.hps_0_f2h_sdram3_data_write                                        (mm_interconnect_1_hps_0_f2h_sdram3_data_write),       //                                                             .write
		.hps_0_f2h_sdram3_data_writedata                                    (mm_interconnect_1_hps_0_f2h_sdram3_data_writedata),   //                                                             .writedata
		.hps_0_f2h_sdram3_data_burstcount                                   (mm_interconnect_1_hps_0_f2h_sdram3_data_burstcount),  //                                                             .burstcount
		.hps_0_f2h_sdram3_data_byteenable                                   (mm_interconnect_1_hps_0_f2h_sdram3_data_byteenable),  //                                                             .byteenable
		.hps_0_f2h_sdram3_data_waitrequest                                  (mm_interconnect_1_hps_0_f2h_sdram3_data_waitrequest)  //                                                             .waitrequest
	);

	cycloneV_soc_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                                      (clk_clk),                                               //                                                    clk_0_clk.clk
		.addVector_0_reset_sink_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                        //                 addVector_0_reset_sink_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                    // hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.addVector_0_avalon_rd1_1_1_1_address                               (addvector_0_avalon_rd1_1_1_1_address),                  //                                 addVector_0_avalon_rd1_1_1_1.address
		.addVector_0_avalon_rd1_1_1_1_waitrequest                           (addvector_0_avalon_rd1_1_1_1_waitrequest),              //                                                             .waitrequest
		.addVector_0_avalon_rd1_1_1_1_burstcount                            (addvector_0_avalon_rd1_1_1_1_burstcount),               //                                                             .burstcount
		.addVector_0_avalon_rd1_1_1_1_read                                  (addvector_0_avalon_rd1_1_1_1_read),                     //                                                             .read
		.addVector_0_avalon_rd1_1_1_1_readdata                              (addvector_0_avalon_rd1_1_1_1_readdata),                 //                                                             .readdata
		.addVector_0_avalon_rd1_1_1_1_readdatavalid                         (addvector_0_avalon_rd1_1_1_1_readdatavalid),            //                                                             .readdatavalid
		.addVector_0_avalon_rd2_address                                     (addvector_0_avalon_rd2_address),                        //                                       addVector_0_avalon_rd2.address
		.addVector_0_avalon_rd2_waitrequest                                 (addvector_0_avalon_rd2_waitrequest),                    //                                                             .waitrequest
		.addVector_0_avalon_rd2_burstcount                                  (addvector_0_avalon_rd2_burstcount),                     //                                                             .burstcount
		.addVector_0_avalon_rd2_read                                        (addvector_0_avalon_rd2_read),                           //                                                             .read
		.addVector_0_avalon_rd2_readdata                                    (addvector_0_avalon_rd2_readdata),                       //                                                             .readdata
		.addVector_0_avalon_rd2_readdatavalid                               (addvector_0_avalon_rd2_readdatavalid),                  //                                                             .readdatavalid
		.addVector_0_avalon_wr_address                                      (addvector_0_avalon_wr_address),                         //                                        addVector_0_avalon_wr.address
		.addVector_0_avalon_wr_waitrequest                                  (addvector_0_avalon_wr_waitrequest),                     //                                                             .waitrequest
		.addVector_0_avalon_wr_write                                        (addvector_0_avalon_wr_write),                           //                                                             .write
		.addVector_0_avalon_wr_writedata                                    (addvector_0_avalon_wr_writedata),                       //                                                             .writedata
		.addVector_1_avalon_rd1_1_1_1_address                               (addvector_1_avalon_rd1_1_1_1_address),                  //                                 addVector_1_avalon_rd1_1_1_1.address
		.addVector_1_avalon_rd1_1_1_1_waitrequest                           (addvector_1_avalon_rd1_1_1_1_waitrequest),              //                                                             .waitrequest
		.addVector_1_avalon_rd1_1_1_1_burstcount                            (addvector_1_avalon_rd1_1_1_1_burstcount),               //                                                             .burstcount
		.addVector_1_avalon_rd1_1_1_1_read                                  (addvector_1_avalon_rd1_1_1_1_read),                     //                                                             .read
		.addVector_1_avalon_rd1_1_1_1_readdata                              (addvector_1_avalon_rd1_1_1_1_readdata),                 //                                                             .readdata
		.addVector_1_avalon_rd1_1_1_1_readdatavalid                         (addvector_1_avalon_rd1_1_1_1_readdatavalid),            //                                                             .readdatavalid
		.addVector_1_avalon_rd2_address                                     (addvector_1_avalon_rd2_address),                        //                                       addVector_1_avalon_rd2.address
		.addVector_1_avalon_rd2_waitrequest                                 (addvector_1_avalon_rd2_waitrequest),                    //                                                             .waitrequest
		.addVector_1_avalon_rd2_burstcount                                  (addvector_1_avalon_rd2_burstcount),                     //                                                             .burstcount
		.addVector_1_avalon_rd2_read                                        (addvector_1_avalon_rd2_read),                           //                                                             .read
		.addVector_1_avalon_rd2_readdata                                    (addvector_1_avalon_rd2_readdata),                       //                                                             .readdata
		.addVector_1_avalon_rd2_readdatavalid                               (addvector_1_avalon_rd2_readdatavalid),                  //                                                             .readdatavalid
		.addVector_1_avalon_wr_address                                      (addvector_1_avalon_wr_address),                         //                                        addVector_1_avalon_wr.address
		.addVector_1_avalon_wr_waitrequest                                  (addvector_1_avalon_wr_waitrequest),                     //                                                             .waitrequest
		.addVector_1_avalon_wr_write                                        (addvector_1_avalon_wr_write),                           //                                                             .write
		.addVector_1_avalon_wr_writedata                                    (addvector_1_avalon_wr_writedata),                       //                                                             .writedata
		.hps_0_f2h_sdram0_data_address                                      (mm_interconnect_2_hps_0_f2h_sdram0_data_address),       //                                        hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                        (mm_interconnect_2_hps_0_f2h_sdram0_data_write),         //                                                             .write
		.hps_0_f2h_sdram0_data_read                                         (mm_interconnect_2_hps_0_f2h_sdram0_data_read),          //                                                             .read
		.hps_0_f2h_sdram0_data_readdata                                     (mm_interconnect_2_hps_0_f2h_sdram0_data_readdata),      //                                                             .readdata
		.hps_0_f2h_sdram0_data_writedata                                    (mm_interconnect_2_hps_0_f2h_sdram0_data_writedata),     //                                                             .writedata
		.hps_0_f2h_sdram0_data_burstcount                                   (mm_interconnect_2_hps_0_f2h_sdram0_data_burstcount),    //                                                             .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                   (mm_interconnect_2_hps_0_f2h_sdram0_data_byteenable),    //                                                             .byteenable
		.hps_0_f2h_sdram0_data_readdatavalid                                (mm_interconnect_2_hps_0_f2h_sdram0_data_readdatavalid), //                                                             .readdatavalid
		.hps_0_f2h_sdram0_data_waitrequest                                  (mm_interconnect_2_hps_0_f2h_sdram0_data_waitrequest)    //                                                             .waitrequest
	);

	cycloneV_soc_mm_interconnect_3 mm_interconnect_3 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                        //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                      //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                       //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                      //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                     //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                      //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                     //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                      //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                     //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                     //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                         //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                       //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                       //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                       //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                      //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                      //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                         //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                       //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                      //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                      //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                        //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                      //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                       //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                      //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                     //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                      //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                     //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                      //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                     //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                     //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                         //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                       //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                       //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                       //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                      //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                      //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                          //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),               // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                   //              onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.onchip_memory2_0_s1_address                                      (mm_interconnect_3_onchip_memory2_0_s1_address),    //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_3_onchip_memory2_0_s1_write),      //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_3_onchip_memory2_0_s1_readdata),   //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_3_onchip_memory2_0_s1_writedata),  //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_3_onchip_memory2_0_s1_byteenable), //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_3_onchip_memory2_0_s1_chipselect), //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_3_onchip_memory2_0_s1_clken)       //                                                           .clken
	);

	cycloneV_soc_mm_interconnect_4 mm_interconnect_4 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                 //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                               //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                               //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                              //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                               //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                              //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                               //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                              //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                              //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                  //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                               //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                               //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                  //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                               //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                               //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                 //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                               //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                               //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                              //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                               //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                              //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                               //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                              //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                              //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                  //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                               //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                               //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                      //                                                     clk_0_clk.clk
		.pll_0_outclk0_clk                                                   (pll_0_outclk0_clk),                                            //                                                 pll_0_outclk0.clk
		.pll_0_outclk1_clk                                                   (pll_0_outclk1_clk),                                            //                                                 pll_0_outclk1.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                           // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.led_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),                               //                               led_reset_reset_bridge_in_reset.reset
		.lwir_ul0304_0_reset_sink_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                           //                lwir_ul0304_0_reset_sink_reset_bridge_in_reset.reset
		.swir_v400_0_reset_sink_reset_bridge_in_reset_reset                  (rst_controller_002_reset_out_reset),                           //                  swir_v400_0_reset_sink_reset_bridge_in_reset.reset
		.addVector_0_slave_1_address                                         (mm_interconnect_4_addvector_0_slave_1_address),                //                                           addVector_0_slave_1.address
		.addVector_0_slave_1_write                                           (mm_interconnect_4_addvector_0_slave_1_write),                  //                                                              .write
		.addVector_0_slave_1_read                                            (mm_interconnect_4_addvector_0_slave_1_read),                   //                                                              .read
		.addVector_0_slave_1_readdata                                        (mm_interconnect_4_addvector_0_slave_1_readdata),               //                                                              .readdata
		.addVector_0_slave_1_writedata                                       (mm_interconnect_4_addvector_0_slave_1_writedata),              //                                                              .writedata
		.addVector_0_slave_1_byteenable                                      (mm_interconnect_4_addvector_0_slave_1_byteenable),             //                                                              .byteenable
		.addVector_0_slave_1_readdatavalid                                   (mm_interconnect_4_addvector_0_slave_1_readdatavalid),          //                                                              .readdatavalid
		.addVector_0_slave_1_waitrequest                                     (mm_interconnect_4_addvector_0_slave_1_waitrequest),            //                                                              .waitrequest
		.addVector_0_slave_1_chipselect                                      (mm_interconnect_4_addvector_0_slave_1_chipselect),             //                                                              .chipselect
		.addVector_1_slave_1_address                                         (mm_interconnect_4_addvector_1_slave_1_address),                //                                           addVector_1_slave_1.address
		.addVector_1_slave_1_write                                           (mm_interconnect_4_addvector_1_slave_1_write),                  //                                                              .write
		.addVector_1_slave_1_read                                            (mm_interconnect_4_addvector_1_slave_1_read),                   //                                                              .read
		.addVector_1_slave_1_readdata                                        (mm_interconnect_4_addvector_1_slave_1_readdata),               //                                                              .readdata
		.addVector_1_slave_1_writedata                                       (mm_interconnect_4_addvector_1_slave_1_writedata),              //                                                              .writedata
		.addVector_1_slave_1_byteenable                                      (mm_interconnect_4_addvector_1_slave_1_byteenable),             //                                                              .byteenable
		.addVector_1_slave_1_readdatavalid                                   (mm_interconnect_4_addvector_1_slave_1_readdatavalid),          //                                                              .readdatavalid
		.addVector_1_slave_1_waitrequest                                     (mm_interconnect_4_addvector_1_slave_1_waitrequest),            //                                                              .waitrequest
		.addVector_1_slave_1_chipselect                                      (mm_interconnect_4_addvector_1_slave_1_chipselect),             //                                                              .chipselect
		.bridge_stSrcMmMaster_0_slave_address                                (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_address),       //                                  bridge_stSrcMmMaster_0_slave.address
		.bridge_stSrcMmMaster_0_slave_write                                  (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_write),         //                                                              .write
		.bridge_stSrcMmMaster_0_slave_read                                   (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_read),          //                                                              .read
		.bridge_stSrcMmMaster_0_slave_readdata                               (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_readdata),      //                                                              .readdata
		.bridge_stSrcMmMaster_0_slave_writedata                              (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_writedata),     //                                                              .writedata
		.bridge_stSrcMmMaster_0_slave_readdatavalid                          (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_readdatavalid), //                                                              .readdatavalid
		.bridge_stSrcMmMaster_0_slave_waitrequest                            (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_waitrequest),   //                                                              .waitrequest
		.bridge_stSrcMmMaster_0_slave_chipselect                             (mm_interconnect_4_bridge_stsrcmmmaster_0_slave_chipselect),    //                                                              .chipselect
		.bridge_stSrcMmMaster_1_slave_address                                (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_address),       //                                  bridge_stSrcMmMaster_1_slave.address
		.bridge_stSrcMmMaster_1_slave_write                                  (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_write),         //                                                              .write
		.bridge_stSrcMmMaster_1_slave_read                                   (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_read),          //                                                              .read
		.bridge_stSrcMmMaster_1_slave_readdata                               (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_readdata),      //                                                              .readdata
		.bridge_stSrcMmMaster_1_slave_writedata                              (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_writedata),     //                                                              .writedata
		.bridge_stSrcMmMaster_1_slave_readdatavalid                          (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_readdatavalid), //                                                              .readdatavalid
		.bridge_stSrcMmMaster_1_slave_waitrequest                            (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_waitrequest),   //                                                              .waitrequest
		.bridge_stSrcMmMaster_1_slave_chipselect                             (mm_interconnect_4_bridge_stsrcmmmaster_1_slave_chipselect),    //                                                              .chipselect
		.led_s1_address                                                      (mm_interconnect_4_led_s1_address),                             //                                                        led_s1.address
		.led_s1_write                                                        (mm_interconnect_4_led_s1_write),                               //                                                              .write
		.led_s1_readdata                                                     (mm_interconnect_4_led_s1_readdata),                            //                                                              .readdata
		.led_s1_writedata                                                    (mm_interconnect_4_led_s1_writedata),                           //                                                              .writedata
		.led_s1_chipselect                                                   (mm_interconnect_4_led_s1_chipselect),                          //                                                              .chipselect
		.lwir_ul0304_0_slave_address                                         (mm_interconnect_4_lwir_ul0304_0_slave_address),                //                                           lwir_ul0304_0_slave.address
		.lwir_ul0304_0_slave_write                                           (mm_interconnect_4_lwir_ul0304_0_slave_write),                  //                                                              .write
		.lwir_ul0304_0_slave_read                                            (mm_interconnect_4_lwir_ul0304_0_slave_read),                   //                                                              .read
		.lwir_ul0304_0_slave_readdata                                        (mm_interconnect_4_lwir_ul0304_0_slave_readdata),               //                                                              .readdata
		.lwir_ul0304_0_slave_writedata                                       (mm_interconnect_4_lwir_ul0304_0_slave_writedata),              //                                                              .writedata
		.lwir_ul0304_0_slave_byteenable                                      (mm_interconnect_4_lwir_ul0304_0_slave_byteenable),             //                                                              .byteenable
		.lwir_ul0304_0_slave_readdatavalid                                   (mm_interconnect_4_lwir_ul0304_0_slave_readdatavalid),          //                                                              .readdatavalid
		.lwir_ul0304_0_slave_waitrequest                                     (mm_interconnect_4_lwir_ul0304_0_slave_waitrequest),            //                                                              .waitrequest
		.lwir_ul0304_0_slave_chipselect                                      (mm_interconnect_4_lwir_ul0304_0_slave_chipselect),             //                                                              .chipselect
		.sw_s1_address                                                       (mm_interconnect_4_sw_s1_address),                              //                                                         sw_s1.address
		.sw_s1_readdata                                                      (mm_interconnect_4_sw_s1_readdata),                             //                                                              .readdata
		.swir_v400_0_slave_address                                           (mm_interconnect_4_swir_v400_0_slave_address),                  //                                             swir_v400_0_slave.address
		.swir_v400_0_slave_write                                             (mm_interconnect_4_swir_v400_0_slave_write),                    //                                                              .write
		.swir_v400_0_slave_read                                              (mm_interconnect_4_swir_v400_0_slave_read),                     //                                                              .read
		.swir_v400_0_slave_readdata                                          (mm_interconnect_4_swir_v400_0_slave_readdata),                 //                                                              .readdata
		.swir_v400_0_slave_writedata                                         (mm_interconnect_4_swir_v400_0_slave_writedata),                //                                                              .writedata
		.swir_v400_0_slave_byteenable                                        (mm_interconnect_4_swir_v400_0_slave_byteenable),               //                                                              .byteenable
		.swir_v400_0_slave_readdatavalid                                     (mm_interconnect_4_swir_v400_0_slave_readdatavalid),            //                                                              .readdatavalid
		.swir_v400_0_slave_waitrequest                                       (mm_interconnect_4_swir_v400_0_slave_waitrequest),              //                                                              .waitrequest
		.swir_v400_0_slave_chipselect                                        (mm_interconnect_4_swir_v400_0_slave_chipselect)                //                                                              .chipselect
	);

	cycloneV_soc_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (0),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_0_outclk1_clk),                     // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (lwir_ul0304_0_st_data),                 //     in_0.data
		.in_0_valid          (lwir_ul0304_0_st_valid),                //         .valid
		.in_0_startofpacket  (lwir_ul0304_0_st_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (lwir_ul0304_0_st_endofpacket),          //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

	cycloneV_soc_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (0),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (pll_0_outclk0_clk),                         // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (swir_v400_0_st_data),                       //     in_0.data
		.in_0_valid          (swir_v400_0_st_valid),                      //         .valid
		.in_0_startofpacket  (swir_v400_0_st_startofpacket),              //         .startofpacket
		.in_0_endofpacket    (swir_v400_0_st_endofpacket),                //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket)    //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk1_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
